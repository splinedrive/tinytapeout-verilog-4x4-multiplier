`timescale 1ns / 1ps
`include "user_module_341493393195532884.v"

module user_module_341493393195532884_tb;

endmodule
